library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity checksum is
    port(
        -- input ports
        i_clk               : in std_logic;
        S_AXIS_T_VALID      : in std_logic;
        S_AXIS_T_LAST       : in std_logic;
        S_AXIS_T_READY      : in std_logic;
        S_AXIS_T_DATA       : in std_logic_vector(7 downto 0);
        i_received_checksum : in std_logic_vector(15 downto 0);
        -- output ports
        o_calc_checksum     : out std_logic_vector(15 downto 0);        
        o_checksum_error    : out std_logic
    );
end checksum;

architecture behavioral of checksum is
type state_type is (EXEC, FINISHED);
signal STATE_REG         : state_type := EXEC; -- por padrão o estado começa como most significant
signal STATE_NEXT        : state_type;

signal CHECK_VALUE_REG     : std_logic_vector(31 downto 0) := (others => '0');
signal CHECK_VALUE_NEXT    : std_logic_vector(31 downto 0) := (others => '0');

signal CHECK_ERROR_REG     : std_logic := '0';
signal CHECK_ERROR_NEXT    : std_logic := '0';

signal CHECK_INTERMED_REG  : std_logic_vector(7 downto 0) := (others => '0');
signal CHECK_INTERMED_NEXT : std_logic_vector(7 downto 0) := (others => '0');

signal CHECK_CALC_REG      : std_logic_vector(31 downto 0) := (others => '0');
signal CHECK_CALC_NEXT     : std_logic_vector(31 downto 0) := (others => '0');

signal CTRL_REG            : std_logic := '0';
signal CTRL_NEXT           : std_logic := '0';

begin
    -- atualização de estado
    clk_process: process(i_clk)
    begin
        if(rising_edge(i_clk)) then
            STATE_REG        <= STATE_NEXT       ;
            CHECK_VALUE_REG    <= CHECK_VALUE_NEXT   ;
            CHECK_ERROR_REG    <= CHECK_ERROR_NEXT   ;
            CHECK_INTERMED_REG <= CHECK_INTERMED_NEXT;
            CHECK_CALC_REG     <= CHECK_CALC_NEXT    ;
            CTRL_REG           <= CTRL_NEXT          ;
        end if;
    end process;

    -- lógica de próximo estado
    next_state: process(STATE_REG, CTRL_REG, S_AXIS_T_VALID, S_AXIS_T_READY, S_AXIS_T_LAST)
    begin
        -- default value
        STATE_NEXT <= STATE_REG;
        CTRL_NEXT    <= CTRL_REG;

        case(STATE_REG) is
            when EXEC =>
                if S_AXIS_T_VALID = '1' and S_AXIS_T_READY = '1' then
                    CTRL_NEXT <= not CTRL_REG;
                    if(S_AXIS_T_LAST = '1') then
                        STATE_NEXT <= FINISHED;
                    end if;
                end if;

            when FINISHED =>
                if S_AXIS_T_VALID = '1' and S_AXIS_T_READY = '1'then
                        STATE_NEXT <= EXEC;
                        CTRL_NEXT <= '1';
                end if;

            when others =>
        end case;
    end process;


    
    datapath: process(STATE_REG,CHECK_VALUE_REG,CHECK_INTERMED_REG, CHECK_CALC_REG, CHECK_ERROR_REG, CTRL_REG, S_AXIS_T_DATA, i_received_checksum, S_AXIS_T_LAST)
    begin
        -- default values
        CHECK_ERROR_NEXT    <= CHECK_ERROR_REG;
        CHECK_INTERMED_NEXT <= CHECK_INTERMED_REG;
        CHECK_VALUE_NEXT    <= CHECK_VALUE_REG;
        CHECK_CALC_NEXT     <= CHECK_CALC_REG;

        case(STATE_REG) is
            when EXEC =>
                if S_AXIS_T_VALID = '1' and S_AXIS_T_READY = '1' and CTRL_REG = '0' then
                    CHECK_INTERMED_NEXT <= S_AXIS_T_DATA;
                    if(S_AXIS_T_LAST = '1') then
                        CHECK_CALC_NEXT <= std_logic_vector(unsigned(CHECK_VALUE_REG)  + unsigned(S_AXIS_T_DATA) - unsigned(i_received_checksum));
                        CHECK_VALUE_NEXT <= std_logic_vector(unsigned(CHECK_VALUE_REG) + unsigned(S_AXIS_T_DATA));
                    end if;
                end if;

                if S_AXIS_T_VALID = '1' and S_AXIS_T_READY = '1' and CTRL_REG = '1' then
                    CHECK_VALUE_NEXT <= std_logic_vector(unsigned(CHECK_VALUE_REG) + unsigned(CHECK_INTERMED_REG & S_AXIS_T_DATA));
                    CHECK_CALC_NEXT  <= std_logic_vector(unsigned(CHECK_VALUE_REG) + unsigned(CHECK_INTERMED_REG & S_AXIS_T_DATA) - unsigned(i_received_checksum));
                end if;
            
            when FINISHED =>
                if((unsigned(CHECK_VALUE_REG) > X"FFFF")) then
                    CHECK_VALUE_NEXT <= std_logic_vector(unsigned(X"0000" & CHECK_VALUE_REG(15 downto 0)) + unsigned(X"0000" & CHECK_VALUE_REG(31 downto 16)));
                    if((unsigned(X"0000" & CHECK_VALUE_REG(15 downto 0)) + unsigned(X"0000" & CHECK_VALUE_REG(31 downto 16))) = X"0000FFFF") then
                        CHECK_ERROR_NEXT <= '0';
                    else
                        CHECK_ERROR_NEXT <= '1';
                    end if;
                else
                    if((unsigned(X"0000" & CHECK_VALUE_REG(15 downto 0))) = X"0000FFFF") then
                        CHECK_ERROR_NEXT <= '0';
                    else
                        CHECK_ERROR_NEXT <= '1';
                    end if;
                end if;

                if((unsigned(CHECK_CALC_REG) > X"FFFF")) then
                    CHECK_CALC_NEXT <= not(std_logic_vector(unsigned(X"0000" & CHECK_CALC_REG(15 downto 0)) + unsigned(X"0000" & CHECK_CALC_REG(31 downto 16))));
                else
                    CHECK_CALC_NEXT <= not(std_logic_vector(unsigned(CHECK_CALC_REG)));
                end if;

                if(S_AXIS_T_LAST = '0') then
                    CHECK_VALUE_NEXT    <= (others => '0');
                    CHECK_ERROR_NEXT    <= '0';
                    CHECK_INTERMED_NEXT <= (others => '0');
                    CHECK_CALC_NEXT     <= (others => '0');
                end if;               
            when others =>
        end case;
    end process;

    o_checksum_error <= CHECK_ERROR_NEXT;
    o_calc_checksum <= CHECK_CALC_NEXT(15 downto 0);

end behavioral;
